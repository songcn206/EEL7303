** Profile: "zenerregulator-Tran"  [ D:\Cadence\SPB_16.6\tools\capture\tclscripts\caplearningresources\hybrid\supportfiles\BasicElectronics\Diode\Designfiles\diode2-pspicefiles\zenerregulator\tran.sim ] 

** Creating circuit file "tran.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
.INC "D:\Cadence\SPB_16.6\tools\capture\tclscripts\caplearningresources\hybrid\supportfiles\BasicElectronics\Diode\Designfiles\diod"
+ "e2-pspicefiles\zenerregulator\tran\tran_profile.inc" 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1m 0 
.STEP LIN PARAM rvariable 1k 10k 2k 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\zenerregulator.net" 


.END
