** Profile: "SCHEMATIC1-AC"  [ D:\OrCAD\bpf\bpf-PSpiceFiles\SCHEMATIC1\AC.sim ] 

** Creating circuit file "AC.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "D:/OrCAD/orcad_10.5_demo/tools/pspice/library/evalaa.lib" 
* From [PSPICE NETLIST] section of D:\OrCAD\OrCAD_10.5_Demo\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 101 1m 1G
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
