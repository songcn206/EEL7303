** Profile: "SCHEMATIC1-zener"  [ D:\CADENCE\SPB_16.5\TOOLS\CAPTURE\FA\Diodes\diode1-PSpiceFiles\SCHEMATIC1\zener.sim ] 

** Creating circuit file "zener.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of D:\Cadence\SPB_16.5\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V1 0 1 0.05 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
