** Profile: "smploscltr-tran80"  [ D:\Cadence\SPB_16.5\tools\capture\FA\OPAmp\opamp-pspicefiles\smploscltr\tran80.sim ] 

** Creating circuit file "tran80.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of D:\Cadence\SPB_16.5\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 50ms 0 1u 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\smploscltr.net" 


.END
