** Profile: "SCHEMATIC1-transient"  [ D:\OrCAD\bpf\bpf-PSpiceFiles\SCHEMATIC1\transient.sim ] 

** Creating circuit file "transient.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "D:/OrCAD/orcad_10.5_demo/tools/pspice/library/evalaa.lib" 
* From [PSPICE NETLIST] section of D:\OrCAD\OrCAD_10.5_Demo\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1 0 1m 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC "..\SCHEMATIC1.net" 


.END
