** Profile: "Diodex-dc"  [ \\pc-alok\d$\public\kit_demo\demo\tools\PSpice\Capture_Samples\paramerized\diodex\diodex-pspicefiles\diodex\dc.sim ] 

** Creating circuit file "dc.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of D:\OrCAD\OrCAD_10.0_Demo\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V1 1 15 0.05 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC "..\Diodex.net" 


.END
